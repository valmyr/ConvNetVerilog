module tb;
parameter SIZE =320, SIZEKer = 5, WIDTH_BIT = 16;
logic clock, nreset,ena,done;
logic signed [WIDTH_BIT-1:0] inpMatrixI          [SIZE-1:0][SIZE-1:0];
logic signed [WIDTH_BIT-1:0] inpMatrixIdinKer    [SIZEKer-1:0][SIZEKer-1:0];

logic signed  [WIDTH_BIT-1:0] convIxKernel ;

logic signed  [WIDTH_BIT-1:0] convIxKernelOut [(SIZE-SIZEKer):0][(SIZE-SIZEKer):0] ;
logic signed  [WIDTH_BIT-1:0] i, j, next,current;
conv2 #(.SIZE(SIZE),.SIZEKer(SIZEKer),.WIDTH_BIT(WIDTH_BIT))top_conv (
    .clock(clock)       ,
    .nreset(nreset)     ,
    .inpMatrixI(inpMatrixI),
    .done(done),
    .convIxKernelOut(convIxKernelOut)
);
initial begin
    $readmemh("simulation/I.txt",inpMatrixI);
    $readmemh("simulation/Kernel.txt",inpMatrixIdinKer);
    clock =0;
    #1nreset = 0;
    #1 nreset = 1;
    do begin 
        #1 clock = ~clock;
    end while(!done);
    $writememh("simulation/IxKernel.txt",convIxKernelOut);
    for(integer i = 0; i < SIZE-SIZEKer+1; i++)begin
        for(integer j = 0; j < SIZE-SIZEKer+1; j++)begin
            $write(convIxKernelOut[i][j]);
        end
        $display("\n");
    end
    for(integer i = 0; i < SIZEKer; i++)begin
        for(integer j = 0; j < SIZEKer; j++)begin
            $write(inpMatrixIdinKer[i][j]);
        end
        $display("\n");
    end
end
endmodule
